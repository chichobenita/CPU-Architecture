---------------------------------------------------------------------------------------------
-- Copyright 2025 Hananya Ribo 
-- Advanced CPU architecture and Hardware Accelerators Lab 361-1-4693 BGU
---------------------------------------------------------------------------------------------
library IEEE;
use ieee.std_logic_1164.all;
USE work.cond_comilation_package.all;



package aux_package is

	component MIPS is
		generic( 
				WORD_GRANULARITY : boolean 	:= G_WORD_GRANULARITY;
				MODELSIM : integer 			:= G_MODELSIM;
				DATA_BUS_WIDTH : integer 	:= 32;
				ITCM_ADDR_WIDTH : integer 	:= G_ADDRWIDTH;
				DTCM_ADDR_WIDTH : integer 	:= G_ADDRWIDTH;
				PC_WIDTH : integer 			:= 10;
				FUNCT_WIDTH : integer 		:= 6;
				DATA_WORDS_NUM : integer 	:= G_DATA_WORDS_NUM;
				CLK_CNT_WIDTH : integer 	:= 16;
				INST_CNT_WIDTH : integer 	:= 16
		);
		PORT(	rst_i		 		:IN		STD_LOGIC;
				clk_i				:IN		STD_LOGIC; 
				BPADDR_i            :IN		STD_LOGIC_VECTOR(7 DOWNTO 0);
				flag_point          :OUT    STD_LOGIC;
			FHCNT_o             :OUT 	STD_LOGIC_VECTOR(7 DOWNTO 0);
			STCNT_o             :OUT	STD_LOGIC_VECTOR(7 DOWNTO 0);
			CLKCNT_o			:OUT	STD_LOGIC_VECTOR(CLK_CNT_WIDTH-1 DOWNTO 0);
			inst_cnt_o 			:OUT	STD_LOGIC_VECTOR(INST_CNT_WIDTH-1 DOWNTO 0);		
			IFpc_o				:OUT    STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
			IFinstruction_o		:OUT    STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			IDpc_o				:OUT    STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
			IDinstruction_o		:OUT    STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			EXpc_o				:OUT    STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
			EXinstruction_o		:OUT    STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			MEMpc_o				:OUT    STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
			MEMinstruction_o	:OUT    STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			WBpc_o				:OUT    STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
			WBinstruction_o		:OUT    STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0)
			
	);		
		
	end component;
---------------------------------------------------------  
	component control is
	PORT( 	
		clk_i 				: IN 	STD_LOGIC;  
		rst_i 				: IN 	STD_LOGIC;
		opcode_i 			: IN 	STD_LOGIC_VECTOR(5 DOWNTO 0);
		RegDst_ctrl_o 		: OUT 	STD_LOGIC_VECTOR(1 DOWNTO 0);
		ALUSrc_ctrl_o 		: OUT 	STD_LOGIC;
		MemtoReg_ctrl_o 	: OUT 	STD_LOGIC;
		RegWrite_ctrl_o 	: OUT 	STD_LOGIC;
		MemRead_ctrl_o 		: OUT 	STD_LOGIC;
		MemWrite_ctrl_o	 	: OUT 	STD_LOGIC;
		Branch_ctrl_o 		: OUT 	STD_LOGIC;
		Bne_ctrl_o 		    : OUT 	STD_LOGIC;
		Beq_ctrl_o 		    : OUT 	STD_LOGIC;
		Jump_ctrl_o         : OUT   STD_LOGIC;
		ALUOp_ctrl_o	 	: OUT 	STD_LOGIC_VECTOR(2 DOWNTO 0)
		);
	end component;
---------------------------------------------------------	
	component dmemory is
		generic(
		DATA_BUS_WIDTH : integer := 32;
		DTCM_ADDR_WIDTH : integer := 8;
		WORDS_NUM : integer := 256
	);
	PORT(	clk_i,rst_i			: IN 	STD_LOGIC;
			dtcm_addr_i 		: IN 	STD_LOGIC_VECTOR(DTCM_ADDR_WIDTH-1 DOWNTO 0);
			dtcm_data_wr_i 		: IN 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			MemRead_ctrl_i  	: IN 	STD_LOGIC;
			MemWrite_ctrl_i 	: IN 	STD_LOGIC;
			dtcm_data_rd_o 		: OUT 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0)
	);
	end component;
---------------------------------------------------------		
	component Execute is
	generic(
		DATA_BUS_WIDTH : integer := 32;
		FUNCT_WIDTH : integer := 6;
		PC_WIDTH : integer := 10
	);
	PORT(	clk_i, rst_i    : IN    STD_LOGIC;
			read_data1_i 	: IN 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			read_data2_i 	: IN 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			sign_extend_i 	: IN 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			funct_i 		: IN 	STD_LOGIC_VECTOR(FUNCT_WIDTH-1 DOWNTO 0);
			ALUOp_ctrl_i 	: IN 	STD_LOGIC_VECTOR(2 DOWNTO 0);
			ALUSrc_ctrl_i 	: IN 	STD_LOGIC;
			pc_plus4_i 		: IN 	STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
			instruction_i 	: IN 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			RegDst_ctrl_i   : IN    STD_LOGIC_VECTOR(1 DOWNTO 0);
			Wr_data_FW_WB_i : IN    STD_LOGIC_VECTOR(31 DOWNTO 0);
			Wr_data_FW_MEM_i: IN    STD_LOGIC_VECTOR(31 DOWNTO 0);
			ForwardA_i      : IN    STD_LOGIC_VECTOR(1 DOWNTO 0);
			ForwardB_i      : IN    STD_LOGIC_VECTOR(1 DOWNTO 0);
			Wr_reg_addr_o   : OUT   STD_LOGIC_VECTOR(4 DOWNTO 0);
			zero_o 			: OUT	STD_LOGIC;
			alu_res_o 		: OUT	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			WriteData_o     : OUT   STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0)
			

	);
	end component;
---------------------------------------------------------		
	component Idecode is
	generic(
		DATA_BUS_WIDTH : integer := 32
	);
	PORT(	clk_i,rst_i		: IN 	STD_LOGIC;
			Stall_ID        : IN    STD_LOGIC;
			instruction_i 	: IN 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			dtcm_data_rd_i 	: IN 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			alu_result_i	: IN 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			RegWrite_ctrl_i : IN 	STD_LOGIC;
			MemtoReg_ctrl_i : IN 	STD_LOGIC;
			JAL_ctrl_i		: IN 	STD_LOGIC;
			pc_plus4_WB_i	: IN 	STD_LOGIC_VECTOR(9 DOWNTO 0);
			--RegDst_ctrl_i 	: IN 	STD_LOGIC_VECTOR(1 DOWNTO 0);
			ForwardA_ID		: IN    STD_LOGIC;
			ForwardB_ID		: IN    STD_LOGIC;
			write_dst_i     : IN 	STD_LOGIC_VECTOR(4 DOWNTO 0);
			Branch_FW_i     : IN    STD_LOGIC_VECTOR(31 DOWNTO 0);
			pc_plus4_i      : IN    STD_LOGIC_VECTOR(9 DOWNTO 0);
			read_data1_o	: OUT 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			read_data2_o	: OUT 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			sign_extend_o 	: OUT 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			Jump_addr_o 	: OUT   STD_LOGIC_VECTOR( 7 DOWNTO 0 );
			PCBranch_addr_o : OUT 	STD_LOGIC_VECTOR(7 DOWNTO 0);
			PCSrc_o		 	: OUT 	STD_LOGIC_VECTOR(1 DOWNTO 0);
			instruction_o 	: OUT 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			write_data_o	: OUT 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0)
		
	);
	end component;
---------------------------------------------------------		
	component Ifetch is
	generic(
		WORD_GRANULARITY : boolean 	:= False;
		DATA_BUS_WIDTH : integer 	:= 32;
		PC_WIDTH : integer 			:= 10;
		NEXT_PC_WIDTH : integer 	:= 8; -- NEXT_PC_WIDTH = PC_WIDTH-2
		ITCM_ADDR_WIDTH : integer 	:= 8;
		WORDS_NUM : integer 		:= 256;
		INST_CNT_WIDTH : integer 	:= 16
	);
	PORT(	
		Stall_IF        : IN    STD_LOGIC;
		clk_i, rst_i 	: IN 	STD_LOGIC;
        Jump_addr_i     : IN    STD_LOGIC_VECTOR(7 DOWNTO 0);
		PCBranch_addr_i : IN    STD_LOGIC_VECTOR(7 DOWNTO 0);
		PCSrc_i		 	: IN 	STD_LOGIC_VECTOR(1 DOWNTO 0);
		pc_o 			: OUT	STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
		pc_plus4_o 		: OUT	STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
		instruction_o 	: OUT	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
		inst_cnt_o 		: OUT	STD_LOGIC_VECTOR(INST_CNT_WIDTH-1 DOWNTO 0)	
	);
	end component;
---------------------------------------------------------
	COMPONENT PLL port(
	    areset		: IN STD_LOGIC  := '0';
		inclk0		: IN STD_LOGIC  := '0';
		c0     		: OUT STD_LOGIC ;
		locked		: OUT STD_LOGIC );
    END COMPONENT;
---------------------------------------------------------	
    COMPONENT shifter is
    generic (
        n           : integer := 32;
        shift_level : integer := 5
    );
    port (
        x    : in std_logic_vector(shift_level-1 downto 0);  -- shift amount
        y    : in std_logic_vector(n-1 downto 0);            -- input vector
        dir  : in std_logic;              -- "0" = SHL, "1" = SHR
        res  : out std_logic_vector(n-1 downto 0)
    );
	END COMPONENT;
---------------------------------------------------------		
	COMPONENT Hazard_forward_Unit IS
	PORT( 
		MemtoReg_EX, MemtoReg_MEM	 		   : IN  STD_LOGIC;
		WriteReg_EX, WriteReg_MEM, WriteReg_WB : IN  STD_LOGIC_VECTOR(4 DOWNTO 0);  -- rt and rd mux output
		RegRs_ID, RegRt_ID 					   : IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		RegRs_EX, RegRt_EX					   : IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		EX_RegWr, MEM_RegWr, WB_RegWr		   : IN  STD_LOGIC;
		BranchBeq_ID, BranchBne_ID			   : IN  STD_LOGIC;
		Stall_IF, Stall_ID, Flush_EX 	 	   : OUT STD_LOGIC;
		ForwardA, ForwardB				       : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		ForwardA_Branch, ForwardB_Branch	   : OUT STD_LOGIC
		);
	END COMPONENT;


end aux_package;

