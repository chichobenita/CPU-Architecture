---------------------------------------------------------------------------------------------
-- Copyright 2025 Hananya Ribo 
-- Advanced CPU architecture and Hardware Accelerators Lab 361-1-4693 BGU
---------------------------------------------------------------------------------------------
-- Ifetch module (provides the PC and instruction 
--memory for the MIPS computer)
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;


ENTITY Ifetch IS
	generic(
		WORD_GRANULARITY : boolean 	:= False;
		DATA_BUS_WIDTH : integer 	:= 32;
		PC_WIDTH : integer 			:= 10;
		NEXT_PC_WIDTH : integer 	:= 8; -- NEXT_PC_WIDTH = PC_WIDTH-2
		ITCM_ADDR_WIDTH : integer 	:= 8;
		WORDS_NUM : integer 		:= 256;
		INST_CNT_WIDTH : integer 	:= 16
	);
	PORT(	
		clk_i, rst_i 	: IN 	STD_LOGIC;
		add_result_i 	: IN 	STD_LOGIC_VECTOR(7 DOWNTO 0);
        Branch_ctrl_i 	: IN 	STD_LOGIC;
		Jump_ctrl_i     : IN    STD_LOGIC;
        zero_i 			: IN 	STD_LOGIC;	
		INT_JMP_MUX_ctrl_i :IN  STD_LOGIC;
		READ_DATA_MEM_i : IN    STD_LOGIC_VECTOR(31 DOWNTO 0);
		TEMP_REG_o      : OUT   STD_LOGIC_VECTOR(31 DOWNTO 0);
		pc_o 			: OUT	STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
		pc_plus4_o 		: OUT	STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
		instruction_o 	: OUT	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
		PC_TO_TEMP_ctrl_i: IN   STD_LOGIC;
		inst_cnt_o 		: OUT	STD_LOGIC_VECTOR(INST_CNT_WIDTH-1 DOWNTO 0)	
	);
END Ifetch;


ARCHITECTURE behavior OF Ifetch IS
	SIGNAL pc_q				  	: STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
	SIGNAL pc_plus4_r 			: STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0);
	SIGNAL itcm_addr_w 			: STD_LOGIC_VECTOR(ITCM_ADDR_WIDTH-1 DOWNTO 0);
	SIGNAL next_pc_w  			: STD_LOGIC_VECTOR(NEXT_PC_WIDTH-1 DOWNTO 0);
	SIGNAL rst_flag_q			: STD_LOGIC;
	SIGNAL inst_cnt_q 			: STD_LOGIC_VECTOR(INST_CNT_WIDTH-1 DOWNTO 0);
	SIGNAL pc_prev_q			: STD_LOGIC_VECTOR(PC_WIDTH-1 DOWNTO 0); 
	SIGNAL jump_addr_w          : STD_LOGIC_VECTOR(NEXT_PC_WIDTH-1 DOWNTO 0);
	SIGNAL next_pc_w1           : STD_LOGIC_VECTOR(NEXT_PC_WIDTH-1 DOWNTO 0);
	SIGNAL INT_JMP_MUX          : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL next_pc_mux  	    : STD_LOGIC_VECTOR(NEXT_PC_WIDTH-1 DOWNTO 0);
	SIGNAL PC_REG_TEMP          : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL sign_extend_PC_TO_TEMP_REG :STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN



--ROM for Instruction Memory
	inst_memory: altsyncram
	GENERIC MAP (
		operation_mode => "ROM",
		width_a => DATA_BUS_WIDTH,
		widthad_a => ITCM_ADDR_WIDTH,
		numwords_a => WORDS_NUM,
		lpm_hint => "ENABLE_RUNTIME_MOD = YES,INSTANCE_NAME = ITCM",
		lpm_type => "altsyncram",
		outdata_reg_a => "UNREGISTERED",
		init_file => "C:\TestPrograms\ModelSim\SW QA - ASM codes\Interrupt based IO\test2\bin\M9K\ITCM.hex",
		intended_device_family => "Cyclone"
	--C:\TestPrograms\ModelSim\SW QA - ASM codes\Interrupt based IO\test2\bin\M9K\ITCM.hex
	)
	PORT MAP (
		clock0     => clk_i,
		address_a  => itcm_addr_w, 
		q_a 	   => instruction_o 
	);
	
	-- Instructions always start on word address - not byte
	pc_q(1 DOWNTO 0) 	<= "00";
	
	-- send address to inst. memory address register
	G1: 
	if (WORD_GRANULARITY = True) generate 		-- i.e. each WORD has unike address
		itcm_addr_w <= next_pc_w;
	elsif (WORD_GRANULARITY = False) generate 	-- i.e. each BYTE has unike address
		itcm_addr_w <= next_pc_w & "00";
	end generate;
		
	-- Adder to increment PC by 4
	pc_plus4_r( 1 DOWNTO 0 )  		 <= "00";
    pc_plus4_r(PC_WIDTH-1 DOWNTO 2)  <= pc_q(PC_WIDTH-1 DOWNTO 2) + 1;
											
	-- Mux to select Branch Address or PC + 4        
	------------------------------------------------------------------------------------				
	next_pc_w1  <= 	(others => '0') WHEN rst_flag_q = '1' ELSE
					add_result_i  	WHEN ((Branch_ctrl_i = '1') AND (
					((zero_i = '1') and (instruction_o(31 DOWNTO 26) = "000100")) or
					((zero_i = '0') and (instruction_o(31 DOWNTO 26) = "000101")))) ELSE
					pc_plus4_r(PC_WIDTH-1 DOWNTO 2);	
					
					
	jump_addr_w <=  (others => '0') WHEN rst_flag_q = '1' ELSE
					instruction_o(7 DOWNTO 0) WHEN instruction_o(31 DOWNTO 26) = "000010" OR instruction_o(31 DOWNTO 26) = "000011" ELSE
					add_result_i WHEN (instruction_o(31 DOWNTO 26) = "000000" AND instruction_o(5 DOWNTO 0) = "001000") ELSE
				    (others => '0');
	next_pc_mux <= next_pc_w1 WHEN (Jump_ctrl_i = '0' and not((instruction_o(31 DOWNTO 26) = "000000" AND instruction_o(5 DOWNTO 0) = "001000"))) ELSE
				    jump_addr_w;
					
	next_pc_w   <=  READ_DATA_MEM_i(9 DOWNTO 2) WHEN  INT_JMP_MUX_ctrl_i = '1' ELSE next_pc_mux;
	-------------------------------------------------------------------------------------
	process (clk_i)
	BEGIN
		IF rising_edge(clk_i) THEN
			rst_flag_q <= rst_i;
		end if;
	end process;
	-------------------------------------------------------------------------------------
	PROCESS (clk_i, rst_i)
	BEGIN
		IF rst_i = '1' THEN
			pc_q(PC_WIDTH-1 DOWNTO 2) <= (OTHERS => '0') ; 
		ELSIF rising_edge(clk_i) THEN
			pc_q(PC_WIDTH-1 DOWNTO 2) <= next_pc_w;	
		END IF;
	END PROCESS;
	
		-- Sign Extend 8-bits to 32-bits
    sign_extend_PC_TO_TEMP_REG <= 	X"000000" & next_pc_w WHEN next_pc_w(7) = '0' ELSE
						X"FFFFFF" & next_pc_w;
	PROCESS (clk_i, rst_i)
	BEGIN
		IF rst_i = '1' THEN
			PC_REG_TEMP <= (OTHERS => '0') ; 
		ELSIF rising_edge(clk_i) THEN
			IF PC_TO_TEMP_ctrl_i = '1' THEN 
			PC_REG_TEMP <= sign_extend_PC_TO_TEMP_REG;	
			END IF;
		END IF;
	END PROCESS;
	
	TEMP_REG_o <= PC_REG_TEMP;
---------------------------------------------------------------------------------------
--						IPC - instruction counter register
---------------------------------------------------------------------------------------
process (clk_i , rst_i)
begin
	if rst_i = '1' then
		pc_prev_q	<=	(others	=> '0');
	elsif falling_edge(clk_i) then
		pc_prev_q	<=	pc_q;
	end if;
end process;
---------------------------------------------------------------------------------------
process (clk_i , rst_i)
begin
	if rst_i = '1' then
		inst_cnt_q	<=	(others	=> '0');
	elsif rising_edge(clk_i) then
		if pc_prev_q = pc_q then
			inst_cnt_q	<=	inst_cnt_q + '1';
		end if;
	end if;
end process;
---------------------------------------------------------------------------------------
	-- copy output signals - allows read inside module
	pc_o 				<= 	pc_q;
	pc_plus4_o 			<= 	pc_plus4_r;
	inst_cnt_o			<=	inst_cnt_q;
END behavior;


